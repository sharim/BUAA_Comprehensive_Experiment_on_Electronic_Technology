module tmp(
	input in,
	output out);

	assign out = ~in;
endmodule // 非门